module RTC_executable(
output [31:0] userTime,
output [31:0] userDate
);

//This module written by getTime.exe

assign userTime=81360;
assign userDate=20323;


endmodule